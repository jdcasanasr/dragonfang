`ifndef RISCV_V_PKG_COMPILED
`define RISCV_V_PKG_COMPILED

package riscv_v_pkg;

	parameter ELEN 			= 64;
	parameter VLEN 			= 64;
	parameter VELEMENTS_MAX = 8;

endpackage

`endif