module tail_encoder
#(
	parameter MASK_LENGTH = 8
)
(
	input 	logic [7:0] mask,
	
	output 	logic [7:0] encoded_mask
);

endmodule 