`ifndef DRAGONFANG_INTEGER_PKG
`define DRAGONFANG_INTEGER_PKG

package dragonfang_integer_pkg;

	// Parameterizable leading bits counter (zero or one).
	`include "C:/Users/jdani/Documents/Thesis/dragonfang/hdl/auxiliary_modules/leading_bits_counter.sv"

endpackage 

`endif